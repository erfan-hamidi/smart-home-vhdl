-- Copyright (C) 2018  Intel Corporation. All rights reserved.
-- Your use of Intel Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Intel Program License 
-- Subscription Agreement, the Intel Quartus Prime License Agreement,
-- the Intel FPGA IP License Agreement, or other applicable license
-- agreement, including, without limitation, that your use is for
-- the sole purpose of programming logic devices manufactured by
-- Intel and sold by Intel or its authorized distributors.  Please
-- refer to the applicable agreement for further details.

-- Generated by Quartus Prime Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition
-- Created on Thu Aug 03 18:46:05 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FinalPorject IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        a : IN STD_LOGIC := '0';
        output1 : OUT STD_LOGIC
    );
END FinalPorject;

ARCHITECTURE BEHAVIOR OF FinalPorject IS
    TYPE type_fstate IS (state1,state2,state3,state4,state5,state7,state8,state9,state10,state11,state6);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,a)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= state1;
            output1 <= '0';
        ELSE
            output1 <= '0';
            CASE fstate IS
                WHEN state1 =>
                    IF ((a = '1')) THEN
                        reg_fstate <= state2;
                    ELSIF (NOT((a = '1'))) THEN
                        reg_fstate <= state1;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state1;
                    END IF;

                    output1 <= '0';
                WHEN state2 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state2;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state2;
                    END IF;

                    output1 <= '0';
                WHEN state3 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state3;
                    END IF;

                    output1 <= '0';
                WHEN state4 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state4;
                    END IF;

                    output1 <= '0';
                WHEN state5 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state3;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state6;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state5;
                    END IF;

                    output1 <= '0';
                WHEN state7 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state8;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state7;
                    END IF;

                    output1 <= '0';
                WHEN state8 =>
                    IF ((a = '1')) THEN
                        reg_fstate <= state5;
                    ELSIF (NOT((a = '1'))) THEN
                        reg_fstate <= state9;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state8;
                    END IF;

                    output1 <= '0';
                WHEN state9 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state10;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state9;
                    END IF;

                    output1 <= '0';
                WHEN state10 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state11;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state5;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state10;
                    END IF;

                    output1 <= '0';
                WHEN state11 =>
                    IF (NOT((a = '1'))) THEN
                        reg_fstate <= state1;
                    ELSIF ((a = '1')) THEN
                        reg_fstate <= state4;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state11;
                    END IF;

                    output1 <= '1';
                WHEN state6 =>
                    IF ((a = '1')) THEN
                        reg_fstate <= state1;
                    ELSIF (NOT((a = '1'))) THEN
                        reg_fstate <= state7;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= state6;
                    END IF;

                    output1 <= '0';
                WHEN OTHERS => 
                    output1 <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
